module test_pipe32;
  reg clk1, clk2;
  integer k;
  pipe_32 pipe_risc32 (clk1, clk2);
  
  initial
    begin
      clk1=0; clk2=0;
      repeat(20) //generate two phase clock
        begin
          #5 clk1=1; #5 clk1=0;
          #5 clk2=1; #5 clk2=0;
        end
    end
  
  initial
    begin
      for(k=0; k<31; k++)
        pipe_32.Reg[k] =k;
      pipe_32.Mem[0] = 32'h2801000a; //ADDI R1, R0, 10
      pipe_32.Mem[1] = 32'h28020014; //ADDI R2, R0, 20
      pipe_32.Mem[2] = 32'h28030019; //ADDI R3, R0, 25
      pipe_32.Mem[3] = 32'h0ce77800; //OR R7, R7, R7 --dummy instruction
      pipe_32.Mem[4] = 32'h0ce77800; //OR R7, R7, R7 --dummy instruction
      pipe_32.Mem[5] = 32'h00222000; //ADD R4, R1, R2
      pipe_32.Mem[6] = 32'h0ce77800; //OR R7, R7, R7 --dummy instruction
      pipe_32.Mem[7] = 32'h00832800; //ADD R5, R4, R3
      pipe_32.Mem[8] = 32'hfc000000; //HLT
      
      pipe_32.HALTED =0;
      pipe_32.PC = 0;
      pipe_32.TAKEN_BRANCH =0;
      #280
      for(k=0; k<6; k++)
        $display("R%1d - %2d",k,pipe_32.Reg[k]);
    end
  
  initial
    begin
      $dumpfile("mips.vcd");
      $dumpvars(0, test_pipe32);
      #300 $finish;
    end
  
      
endmodule
